library verilog;
use verilog.vl_types.all;
entity memory is
    port(
        clock           : in     vl_logic;
        sram_1_addressline_1: in     vl_logic_vector(8 downto 0);
        sram_1_addressline_2: in     vl_logic_vector(8 downto 0);
        sram_2_addressline_1: in     vl_logic_vector(8 downto 0);
        sram_2_addressline_2: in     vl_logic_vector(8 downto 0);
        sram_3_addressline_1: in     vl_logic_vector(8 downto 0);
        sram_3_addressline_2: in     vl_logic_vector(8 downto 0);
        sram_4_addressline_1: in     vl_logic_vector(8 downto 0);
        sram_4_addressline_2: in     vl_logic_vector(8 downto 0);
        sram_1_readline_1: out    vl_logic_vector(47 downto 0);
        sram_1_readline_2: out    vl_logic_vector(47 downto 0);
        sram_2_readline_1: out    vl_logic_vector(47 downto 0);
        sram_2_readline_2: out    vl_logic_vector(47 downto 0);
        sram_3_readline_1: out    vl_logic_vector(47 downto 0);
        sram_3_readline_2: out    vl_logic_vector(47 downto 0);
        sram_4_readline_1: out    vl_logic_vector(47 downto 0);
        sram_4_readline_2: out    vl_logic_vector(47 downto 0);
        sram1_WriteAddress1: in     vl_logic_vector(8 downto 0);
        sram1_WriteAdress2: in     vl_logic_vector(8 downto 0);
        sram2_WriteAddress1: in     vl_logic_vector(8 downto 0);
        sram2_WriteAdress2: in     vl_logic_vector(8 downto 0);
        sram3_WriteAddress1: in     vl_logic_vector(8 downto 0);
        sram3_WriteAdress2: in     vl_logic_vector(8 downto 0);
        sram4_WriteAddress1: in     vl_logic_vector(8 downto 0);
        sram4_WriteAdress2: in     vl_logic_vector(8 downto 0);
        sram1_WriteBus1 : out    vl_logic_vector(47 downto 0);
        sram1_WriteBus2 : out    vl_logic_vector(47 downto 0);
        sram2_WriteBus1 : out    vl_logic_vector(47 downto 0);
        sram2_WriteBus2 : out    vl_logic_vector(47 downto 0);
        sram3_WriteBus1 : out    vl_logic_vector(47 downto 0);
        sram3_WriteBus2 : out    vl_logic_vector(47 downto 0);
        sram4_WriteBus1 : out    vl_logic_vector(47 downto 0);
        sram4_WriteBus2 : out    vl_logic_vector(47 downto 0);
        yram_WriteAddress: in     vl_logic_vector(10 downto 0);
        Y_addressline_1 : in     vl_logic_vector(10 downto 0);
        ReadAddress2    : in     vl_logic_vector(10 downto 0);
        ReadBus2        : out    vl_logic_vector(255 downto 0);
        ReadBus1        : out    vl_logic_vector(255 downto 0);
        y_WriteBus      : in     vl_logic_vector(255 downto 0);
        WE_1            : in     vl_logic;
        WE_2            : in     vl_logic;
        WE_3            : in     vl_logic;
        WE_4            : in     vl_logic;
        WE_Y            : in     vl_logic;
        WE_I            : in     vl_logic;
        WriteAddress_I  : in     vl_logic_vector(7 downto 0);
        I_sram_addressline_1: in     vl_logic_vector(7 downto 0);
        I_sram_ReadAddress2: in     vl_logic_vector(7 downto 0);
        I_WriteBus      : in     vl_logic_vector(191 downto 0);
        I_sram_ReadBus2 : out    vl_logic_vector(191 downto 0);
        I_sram_ReadBus1 : out    vl_logic_vector(191 downto 0)
    );
end memory;
